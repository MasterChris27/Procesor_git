----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    15:18:45 05/15/2018 
-- Design Name: 
-- Module Name:    IO - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity IO is
    Port ( Clk : in  STD_LOGIC;
			  Bus_control : in std_logic_vector(1 downto 0);
           Bus_data : in  STD_LOGIC_VECTOR (15 downto 0);
           Bus_address : in  STD_LOGIC_VECTOR (15 downto 0));
end IO;

architecture Behavioral of IO is

begin


end Behavioral;

